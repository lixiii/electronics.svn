* Version 1.67 Copyright ? Linear Technology Corp. 5/19/04. All rights reserved. [Spice2]
* Node List: IN+(3) IN-(2) VCC(7) VEE(4) OUT(6)
.SUBCKT LT6220 3 2 7 4 6
CCM1 162 0 0.001
CG2 158 0 1n
CG3 159 0 5e-7
CG5 164 0 1.26582e-8
CG7 165 0 1e-10
CIN1 3 2 0.1f
CIN2 0 3 2p
CIN3 2 0 2p
CPSN 179 0 10p
CPSN2 178 0 1e-6
CPSP 181 0 10p
CPSP2 180 0 1e-6
CVM 175 0 1E5
DIN1 108 7 DIODE
DIN2 103 7 DIODE
DIN3 4 108 DIODE
DIN4 4 103 DIODE
DIN5 103 108 DIODE
DIN6 108 103 DIODE
DVLIM1 177 144 DVLIM
DVLIM2 145 177 DVLIM
DVNF 146 0 DVNOI
DVNFX 147 0 DVNOIX
EICM1 153 0 2 0 1
EICM2 154 0 3 0 1
EILIM1 125 122 177 155 1E5
EILIM2 124 120 177 155 -1E5
EIN1 106 0 105 0 1
EIN2 104 0 103 0 1
EPWR1 135 0 177 155 1E5
EPWR2 136 0 177 155 1E5
ESRLIM1 141 143 103 105 0
ESRLIM2 140 142 105 103 0
ESRLIM3 140 138 157 156 499.091
ESRLIM4 141 139 156 157 499.091
EVCC 161 0 7 0 1
EVEE 167 0 4 0 1
EVNOI1 107 108 0 148 1
EVNOI2 109 107 146 147 1
FVLIM1 177 0 VVLIM1 -1E7
FVLIM2 177 0 VVLIM2 1E7
GCM2 0 163 170 175 0.000446684
GCM3 0 162 163 0 6.2832
GCMO1 0 159 162 0 6.2832
GG2 0 158 157 156 0.313589
GG3 0 159 158 0 10
GG5 0 164 159 0 6.2832
GG7 0 165 164 0 6.2832
GILIM 158 0 128 0 0.01
GINOI1 103 0 0 129 1m
GINOI2 110 0 0 130 1m
GOUT2 0 177 169 0 10
GPSN2 0 179 4 175 0.000794328
GPSN4 0 178 179 0 6.2832
GPSNO2 0 177 178 0 10
GPSP2 0 181 7 175 0.000794328
GPSP4 0 180 181 0 6.2832
GPSPO2 0 177 180 0 10
GPWR1 133 0 177 155 100
GPWR2 134 0 177 155 100
GSHD3 4 7 119 0 1
GZP1 167 168 165 0 0.1
GZP3 167 169 168 0 0.1
HIN1 113 156 VIN1 100
HIN2 118 157 VIN2 100
HIN3 116 117 VIN3 100
HIN4 112 115 VIN4 100
IBIAS1 105 0 1.5e-8
IBIAS2 103 0 1.5e-8
IDUM1 148 0 0
IDUM2 130 129 0
IPWR 7 4 0.001
ISLEW 111 0 10mA
IVNF 0 146 1A
IVNFX 0 147 1A
LCM2 127 0 0.00530516
LCMX 126 163 100
LPSN2 131 0 1.59155e-8
LPSP2 132 0 1.59155e-8
LZP2 149 167 2.27205e-7
LZP4 150 167 1.76839e-11
Q1 156 106 116 0 NPN1
Q2 157 104 112 0 NPN1
RCM2 163 127 1k
RCM3 162 0 0.159155
RCMX 126 0 0.1
RCMX2 163 126 1E8
RG2 158 0 159155
RG3 159 0 0.159155
RG5 164 0 0.159155
RG7 165 0 0.159155
RICM1 153 170 1k
RICM2 154 170 1k
RILIM 128 0 1
RIN1 108 3 0.1
RIN2 103 2 0.1
RINOI1 129 0 38.6473
RINOI2 130 0 38.6473
ROUT2 177 0 0.1
ROUT3 176 155 0.01
RPSN2 179 131 1k
RPSN22 131 0 1E8
RPSN4 178 0 0.159155
RPSP2 181 132 1k
RPSP22 132 0 1E8
RPSP4 180 0 0.159155
RPWR1 133 161 1E6
RPWR2 134 167 1E6
RSENSE 155 177 0.01
RSHD1 119 0 1
RVH1 161 175 1k
RVH2 175 167 1k
RVNOI 0 148 6038.45
RZP1 168 149 10
RZP4 149 167 14275.7
RZP5 169 150 10
RZP8 150 167 1.11111
SHD2 137 119 7 4 SHDN2X
SHD8 152 6 7 4 SHDNO2
SILIM1 128 123 122 0 SILIM
SILIM2 128 121 120 0 SILIM
SPWR1 7 133 135 0 SPWR
SPWR2 4 134 136 0 SPWRX
SSRLIM1 156 157 138 0 SSRLIM
SSRLIM2 156 157 139 0 SSRLIM
VILIM1 125 0 35
VILIM2 124 0 35
VILIM3 123 0 10000
VILIM4 121 0 -10000
VIN1 114 113 0
VIN2 114 118 0
VIN3 117 111 0
VIN4 115 111 0
VINPUT 114 0 100
VNF 109 110 83.3788uV
VOS 105 110 200u
VSHD7 152 176 0
VSHDN 137 0 0.000999
VSRLIM1 142 0 20
VSRLIM2 143 0 20
VVLIM1 161 144 1.2535
VVLIM2 145 167 1.2235
.MODEL NPN1 NPN(BF=1E11 BR=1E11 AF=0 KF=0 XTI=0 CJC=1f CJE=1f CJS=1f )
.MODEL SHDN VSWITCH(ROFF=1E7 RON=0.001 VON=1.80V VOFF=2.00V)
.MODEL SHDNX VSWITCH(ROFF=1E7 RON=0.001 VON=2.00V VOFF=1.80V)
.MODEL SHDNO VSWITCH(ROFF=1000000.00 RON=0.001 VON=1.80V VOFF=2.00V)
.MODEL SHDNO2 VSWITCH(ROFF=1000000.00 RON=0.001 VON=1.10V VOFF=0.90V)
.MODEL SHDNOX VSWITCH(ROFF=1000000.00 RON=0.001 VON=2.00V VOFF=1.80V)
.MODEL SHDN2 VSWITCH(ROFF=1E7 RON=0.001 VON=1.10V VOFF=0.90V)
.MODEL SHDN2X VSWITCH(ROFF=1E7 RON=0.001 VON=0.90V VOFF=1.10V)
.MODEL SBIAS VSWITCH(ROFF=1E7 RON=0.001 VON=0.80V VOFF=1.00V)
.MODEL SBIAS2 VSWITCH(ROFF=1E7 RON=0.001 VON=1.00V VOFF=0.80V)
.MODEL SBIASX VSWITCH(ROFF=1E7 RON=0.001 VON=1.00V VOFF=0.80V)
.MODEL SBIAS2X VSWITCH(ROFF=1E7 RON=0.001 VON=0.80V VOFF=1.00V)
.MODEL SSRLIM VSWITCH(ROFF=1E7 RON=0.01 VON=-0.1 VOFF=0.5)
.MODEL SILIM VSWITCH(ROFF=1E7 RON=0.001 VON=-3V VOFF=0.4V)
.MODEL SPWR VSWITCH(ROFF=1G RON=0.1 VON=12V VOFF=-12V)
.MODEL SPWRX VSWITCH(ROFF=1G RON=0.1 VON=-12V VOFF=12V)
.MODEL DIODE D(KF=0 RS=0)
.MODEL DVLIM D(IS=1E-24 KF=0 RS=0 XTI=0)
.MODEL DVNOIX D(KF=0 RS=0)
.MODEL DIDEAL D(KF=0 RS=0 XTI=0)
.MODEL DVNOI D(RS=0 KF= 1.49279e-11)
.ENDS LT6220